module LCD_interface(
    input logic clk, rstN,
    input logic 
)