module master 
(
    input logic clk, rstN,
    output logic control,write_data,valid,last,
    input logic read_data, ready
);


endmodule: master