bus_state