module interconnect #(
    parameters
) (
    //arbiter
    input Master,
    input Slave, 
    
);
    
endmodule