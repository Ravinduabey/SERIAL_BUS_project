module arbiter(
    input logic clk,
	 input logic rstn,
    input logic m1_in,
	 input logic m2_in,
	 output logic m1_out,
	 output logic m2_out,
	 input logic ready,
	 output logic buscontrol
);



endmodule : arbiter